pBAV       4  ��   @  ����n.@   ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  .    ��������  n@$ $$      �����_   � � � �   @% %%      �����S   � � � �   Z@+ &&      �����_   � � � �   n@; ''      �����_   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �   ~ @"                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       