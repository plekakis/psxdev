pBAV       p� �� _  @  ����P �@   ��������P �@   ��������P �@   ��������P �@   ��������P �@   ��������P �@   ��������P �@   ��������P �@   ��������P �@   ��������P �@   ��������P �@   ��������P �@   ��������P �@   ��������P �@   �������� �@   ��������	 �@   ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������  $  +    �����	   � � � �   -0 *7    �����	   � � � �   << 6C    �����	   � � � �   KH BO    �����	   � � � �   ZT N    �����	   � � � �             ��        � � � �             ��        � � � �             ��        � � � �             ��        � � � �             ��        � � � �             ��        � � � �             ��        � � � �             ��        � � � �             ��        � � � �             ��        � � � �             ��        � � � �   $  +    �����	  � � � �   -0 *7    �����	  � � � �   << 6C    �����	  � � � �   KH BO    �����	  � � � �   ZT N    �����	  � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �   $  +    �����	  � � � �   -0 *7    �����	  � � � �   << 6C    �����	  � � � �   KH BO    �����	  � � � �   ZT N    �����	  � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �   $  +    �����	  � � � �   -0 *7    �����	  � � � �   << 6C    �����	  � � � �   KH BO    �����	  � � � �   ZT N    �����	  � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �   $  +    �����	  � � � �   -0 *7    �����	  � � � �   << 6C    �����	  � � � �   KH BO    �����	  � � � �   ZT N    �����	  � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �   $  +    �����	  � � � �   -0 *7    �����	  � � � �   << 6C    �����	  � � � �   KH BO    �����	  � � � �   ZT N    �����	  � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �   $  +    �����	  � � � �   -0 *7    �����	  � � � �   << 6C    �����	  � � � �   KH BO    �����	  � � � �   ZT N    �����	  � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �   $  +    �����	  � � � �   -0 *7    �����	  � � � �   << 6C    �����	  � � � �   KH BO    �����	  � � � �   ZT N    �����	  � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �   $  +    �����	  � � � �   -0 *7    �����	  � � � �   << 6C    �����	  � � � �   KH BO    �����	  � � � �   ZT N    �����	  � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �   $  +    �����		  � � � �   -0 *7    �����		  � � � �   << 6C    �����		  � � � �   KH BO    �����		  � � � �   ZT N    �����		  � � � �             ��    	   � � � �             ��    	   � � � �             ��    	   � � � �             ��    	   � � � �             ��    	   � � � �             ��    	   � � � �             ��    	   � � � �             ��    	   � � � �             ��    	   � � � �             ��    	   � � � �             ��    	   � � � �   $  +    �����	
  � � � �   -0 *7    �����	
  � � � �   << 6C    �����	
  � � � �   KH BO    �����	
  � � � �   ZT N    �����	
  � � � �             ��    
   � � � �             ��    
   � � � �             ��    
   � � � �             ��    
   � � � �             ��    
   � � � �             ��    
   � � � �             ��    
   � � � �             ��    
   � � � �             ��    
   � � � �             ��    
   � � � �             ��    
   � � � �   $  +    �����	  � � � �   -0 *7    �����	  � � � �   << 6C    �����	  � � � �   KH BO    �����	  � � � �   ZT N    �����	  � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �   $  +    �����	  � � � �   -0 *7    �����	  � � � �   << 6C    �����	  � � � �   KH BO    �����	  � � � �   ZT N    �����	  � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �   $  +    �����	  � � � �   -0 *7    �����	  � � � �   << 6C    �����	  � � � �   KH BO    �����	  � � � �   ZT N    �����	  � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �   @$ !%    ��� � 	 � � � �   @& &'    ��� M 
 � � � �   6' '(    ��� �  � � � �   "= )*    ��� �  � � � �   :5 -.    ��� �  � � � �   R3 01    ��� �  � � � �   ^2 23    ��� �  � � � �   T* 45    ��� �  � � � �   T. ./    ��� �  � � � �   T1 12    ��� �  � � � �   TA AB    ��� �  � � � �   '8 89    ��� �  � � � �   'C CD    ��� �  � � � �   Z% %&    ��� �  � � � �   T7 78    ��� �  � � � �   ZcH HP    ��� �  � � � �   {      ��� �_  � � � �   n     ��� �  � � � �           ��� �  � � � �   " !"    ��� �  � � � �   20 #$    ���*M  � � � �   2a2 %'    ���*M  � � � �   @( ((    ��� �_  � � � �   @* )+    ��� �_  � � � �   @, ,-    ��� �_  � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �             ��       � � � �   �.�& 	�*0.`�|T ���
��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                