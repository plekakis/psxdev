pBAV       `w ��   @  ����@@   ��������,@@   ��������<@@   ��������0@   ��������4@d   ��������*@P   ��������&@@   ��������*@@   ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  R@& $$      ������   � � � �   N@& &&      ������   � � � �   X, **      ��!���   � � � �   <X0 ..      ������   � � � �   d,5 11      ��w�	�   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �   @6�     ��Հh�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @;        ���)�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @4        �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @+        ������  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @?a       ������ 	 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @B6       ������ 
 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @Hy       ����f�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   tj�� 8�HfD�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        