pBAV       @� ��   @  ����R�D*   ��������\�D@   ��������\�DV   ��������X�DH   ��������R�D@   ��������R�DH   ��������P�D@   ��������\�D:   ��������X�DP   ��������R�D@   ��������P�D    ��������P�Dd   ��������P�D4   ��������L�D$   ��������P�D0   ��������n�D@   ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    ��������  �D    �������� \@TE    �����_   � � � �  \@H6D    �����_   � � � �  \@< 5    �����_   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  Z@TE    �����_  � � � �  Z@H 6D    �����_  � � � �  Z@< 5    �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  Z@U{E    �����_  � � � �  Z@Is6D    �����_  � � � �  Z@={ 5    �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  d@R       ����KQ  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  d@<     ����IR  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  d@D~     ����IQ  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  Z@FW       ����JQ  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  d@@       �����P  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  d@F       �����Q 	 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  x@<      �����P	 
 � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �  d@E        �����_
  � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �  t@C        ��w��O  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@Et       ����IQ  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@<        ����P  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  t@< <<      �����_  � � � �  t@>:>>      �����_  � � � �  V@_ @@    �����_  � � � �  V@` AA    �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  DNH@HH      ��Ԁ@  � � � �  DNJ JJ      ��Ԁ@  � � � �  H<  .      �����O  � � � �  H ; ;;      ��	�	L  � � � �  > < <<      ��X�	P  � � � �  > > >>      ��W�	P  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    ���� 
~��6 @� 4�\�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          