pBAV       �� ��   @  ����w�@   ��������w�@   ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  w�    ��������  @$ !%    �����   � � � �   @& &&    �����   � � � �   6' '(    �����   � � � �   "= )*    �����   � � � �   :5 --    �����   � � � �   R3 00    �����   � � � �   ^2 22    �����   � � � �   T* 44    �����   � � � �   T. ..    �����   � � � �   T1 11    �����  
 � � � �   TA AA    �����   � � � �   '8 88    �����   � � � �   'C CC    �����   � � � �   Z% %%    �����   � � � �   T7 77    �����   � � � �   ZcH HJ    �����_   � � � �   {      ��� �  � � � �   n(     ��� �  � � � �      !    ��� �  � � � �   " !#    ��� �  � � � �   20 #%    ���*M  � � � �   2a2 %'    ���*M  � � � �   @( ()    ��� �  � � � �   @* )+    ��� M  � � � �   @, ,-    ��� �  � � � �  @<  x<  �����_ 	 � � � �   @<  x    �����_ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   $ 0.`�|T$ ���
��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          