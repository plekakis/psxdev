pBAV       �  ��   @  ����n@@   ��������n@@   ��������n@@   ��������n@    ��������n@@   ��������n@   ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    ��������  @    �������� F@Dz     ����)Q   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  d@T        �����N  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  d@<        �����Q  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  d@<       �����Q  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  d@<       �����Q  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  d@<       �����Q  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   �� Bf                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      