pBAV       �o ��   @  ����d�@   ��������d�@   ��������n�@   ��������d�@   ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  n@$ $$      ������   � � � �   n@* **      ��"�i�   � � � �  n@> 22      ������   � � � �  d@9 33      ������   � � � �  d@; 44      ������   � � � �  x@8 11      ������   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  n@<  <      �����_  � � � �  i@H =H      �����_ 	 � � � �  d@T I      �����_ 
 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  p@<  5      ������  � � � �  k@< 6C      ������  � � � �  h@< DJ      ������  � � � �  a@< KO      ������  � � � �  Z@< PT      ������  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   n@0        ������  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   �� r� X�X��  
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        